// https://www.edaplayground.com/x/iDDu

module negedge_3bit_up_counter_test();
    reg CLK, not_RST, not_PRE;
    wire Q0, Q1, Q2;

    negedge_3bit_up_counter negedge_3bit_up_counter_dut(CLK, not_RST, not_PRE, Q0, Q1, Q2);

    initial begin
        CLK = 1;
        forever #5 CLK = ~CLK;
    end
    initial begin
        not_RST = 0; not_PRE = 1; #10;
        not_RST = 1; not_PRE = 1; #80;
        $finish;
    end
    initial begin
        $dumpfile("test.vcd");
        $dumpvars(1, negedge_3bit_up_counter_test);
    end
endmodule
